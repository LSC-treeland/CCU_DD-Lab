module add(a, b, c, d, res);

	input [3:0] a, b ,c ,d;	
	output [5:0] res;	
	assign res = a + b + c + d;	

endmodule

